*Automatic generated instance fron ../../tech/scripts/genxdut dig
adut [clk
+ cmp
+ ]
+ [b.4
+ b.3
+ b.2
+ b.1
+ b.0
+ reset
+ ] null dut
.model dut d_cosim simulation="../dig.so" delay=10p

* Inputs
Rsvi0 clk 0 1G
Rsvi1 cmp 0 1G

* Outputs
Rsvi2 b.4 0 1G
Rsvi3 b.3 0 1G
Rsvi4 b.2 0 1G
Rsvi5 b.1 0 1G
Rsvi6 b.0 0 1G
Rsvi7 reset 0 1G

E_STATE_b dec_b 0 value={( 0 
+ + 16*v(b.4)/AVDD
+ + 8*v(b.3)/AVDD
+ + 4*v(b.2)/AVDD
+ + 2*v(b.1)/AVDD
+ + 1*v(b.0)/AVDD
+)/1000}
.save v(dec_b)

.save v(reset)

