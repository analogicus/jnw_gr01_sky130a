magic
tech sky130A
magscale 1 2
timestamp 1744207573
<< viali >>
rect -41 10799 33 10873
rect 7 8365 85 8443
rect 1736 8240 1928 8367
rect 364 7714 604 7842
rect 3868 7602 4108 7830
rect 4354 6437 4431 6514
rect 4356 4290 4456 4402
rect 342 3938 570 4166
rect 3848 3898 4088 4032
rect 5100 3028 5200 3128
rect 5111 1877 5194 1960
rect 6987 1709 7053 1775
rect -24 632 65 721
rect 5136 634 5221 719
rect 6930 540 7026 636
<< metal1 >>
rect -47 10879 39 10885
rect -47 10787 39 10793
rect 290 10752 296 10920
rect 382 10752 388 10920
rect 312 10322 480 10328
rect 124 10192 130 10284
rect 222 10192 228 10284
rect 312 10194 480 10200
rect 672 9618 864 10330
rect 1606 9618 1798 9620
rect 672 9316 1798 9618
rect 154 8936 160 9000
rect 224 8936 230 9000
rect 672 8824 864 9316
rect 2370 9134 2376 9326
rect 2536 9134 2568 9326
rect 2120 9040 2288 9046
rect 2120 8866 2288 8872
rect 2376 8828 2568 9134
rect 672 8720 864 8766
rect 1 8449 91 8455
rect 1 8353 91 8359
rect 300 8320 306 8488
rect 396 8450 402 8488
rect 396 8320 442 8450
rect 1992 8384 2056 8390
rect 351 8258 442 8320
rect 1724 8367 1940 8373
rect 351 8252 554 8258
rect 1724 8252 1736 8367
rect 351 8240 1736 8252
rect 1928 8252 1940 8367
rect 1992 8314 2056 8320
rect 1928 8251 3172 8252
rect 4247 8251 4253 8301
rect 1928 8240 4253 8251
rect 351 8182 4253 8240
rect 351 8180 3172 8182
rect 351 8171 554 8180
rect 414 7848 554 8171
rect 1763 8157 1902 8180
rect 4247 8179 4253 8182
rect 4375 8251 4381 8301
rect 4375 8182 5734 8251
rect 4375 8179 4381 8182
rect 352 7842 616 7848
rect 352 7714 364 7842
rect 604 7714 616 7842
rect 352 7708 616 7714
rect 3856 7830 4120 7836
rect 3856 7602 3868 7830
rect 4108 7602 4120 7830
rect 3856 7596 4120 7602
rect 3868 6330 4108 7596
rect 5665 6707 5734 8182
rect 4730 6520 4842 6524
rect 5361 6520 5877 6707
rect 4342 6514 5877 6520
rect 4342 6437 4354 6514
rect 4431 6437 5877 6514
rect 4342 6431 5877 6437
rect 336 6090 4108 6330
rect 336 4166 576 6090
rect 4730 4514 4842 6431
rect 5361 6243 5877 6431
rect 5469 6237 5877 6243
rect 4350 4402 4462 4414
rect 4730 4402 5632 4514
rect 4350 4290 4356 4402
rect 4456 4346 5632 4402
rect 4456 4290 4842 4346
rect 4350 4278 4462 4290
rect 336 3938 342 4166
rect 570 3938 576 4166
rect 336 3926 576 3938
rect 3836 4032 4100 4038
rect 3836 3898 3848 4032
rect 4088 3898 4100 4032
rect 3836 3892 4100 3898
rect 3895 3668 4041 3892
rect -30 727 71 733
rect -30 620 71 626
rect 282 592 288 760
rect 389 592 395 760
rect 3883 710 4094 3668
rect 5464 3576 5632 4346
rect 5464 3408 7464 3576
rect 5464 3162 5632 3408
rect 5094 3134 5206 3140
rect 5094 3016 5206 3022
rect 5434 2994 5440 3162
rect 5552 2994 5632 3162
rect 5302 2468 5308 2532
rect 5372 2468 5378 2532
rect 5105 1966 5200 1972
rect 5105 1865 5200 1871
rect 5434 1822 5440 2014
rect 5535 1822 5541 2014
rect 5824 1894 6016 2594
rect 6102 2108 6108 2172
rect 6172 2108 7208 2172
rect 6981 1781 7059 1787
rect 7144 1762 7208 2108
rect 7296 1826 7464 3408
rect 6981 1697 7059 1703
rect 7266 1658 7272 1826
rect 7350 1658 7464 1826
rect 5320 1442 5384 1448
rect 5314 1438 5384 1442
rect 5312 1413 5384 1438
rect 5312 1378 5390 1413
rect 4730 1174 4938 1228
rect 5312 1174 5384 1378
rect 4730 1102 5384 1174
rect 4730 1040 4938 1102
rect 4732 1038 4938 1040
rect 5444 1072 5636 1490
rect 7138 1126 7144 1190
rect 7208 1126 7214 1190
rect 5444 880 6016 1072
rect 5824 760 6016 880
rect 5130 725 5227 731
rect 769 630 4094 710
rect 769 578 2695 630
rect 2747 578 4094 630
rect 5124 628 5130 725
rect 5227 628 5233 725
rect 5130 622 5227 628
rect 5434 592 5440 760
rect 5537 592 5543 760
rect 769 499 4094 578
rect 5824 568 5927 760
rect 6016 568 6022 760
rect 6924 642 7032 648
rect 6924 528 7032 534
rect 7266 492 7272 684
rect 7380 492 7386 684
rect 7656 532 7848 1248
rect 166 182 172 246
rect 224 182 230 246
rect 5326 241 5378 247
rect 296 -4 464 208
rect 5326 183 5378 189
rect 2646 -4 3098 164
rect 296 -10 3098 -4
rect 5450 -10 5618 208
rect 6577 114 6782 248
rect 6577 50 7208 114
rect 6577 23 6782 50
rect 6580 20 6782 23
rect 296 -81 5618 -10
rect 296 -133 1991 -81
rect 2065 -133 5618 -81
rect 296 -172 5618 -133
rect 2652 -178 5618 -172
<< via1 >>
rect -47 10873 39 10879
rect -47 10799 -41 10873
rect -41 10799 33 10873
rect 33 10799 39 10873
rect -47 10793 39 10799
rect 296 10752 382 10920
rect 130 10192 222 10284
rect 312 10200 480 10322
rect 160 8936 224 9000
rect 2376 9134 2536 9326
rect 2120 8872 2288 9040
rect 672 8766 864 8824
rect 1 8443 91 8449
rect 1 8365 7 8443
rect 7 8365 85 8443
rect 85 8365 91 8443
rect 1 8359 91 8365
rect 306 8320 396 8488
rect 1992 8320 2056 8384
rect 4253 8179 4375 8301
rect 3978 3906 4042 3970
rect -30 721 71 727
rect -30 632 -24 721
rect -24 632 65 721
rect 65 632 71 721
rect -30 626 71 632
rect 288 592 389 760
rect 5094 3128 5206 3134
rect 5094 3028 5100 3128
rect 5100 3028 5200 3128
rect 5200 3028 5206 3128
rect 5094 3022 5206 3028
rect 5440 2994 5552 3162
rect 5308 2468 5372 2532
rect 5105 1960 5200 1966
rect 5105 1877 5111 1960
rect 5111 1877 5194 1960
rect 5194 1877 5200 1960
rect 5105 1871 5200 1877
rect 5440 1822 5535 2014
rect 6108 2108 6172 2172
rect 6981 1775 7059 1781
rect 6981 1709 6987 1775
rect 6987 1709 7053 1775
rect 7053 1709 7059 1775
rect 6981 1703 7059 1709
rect 7272 1658 7350 1826
rect 2695 578 2747 630
rect 5130 719 5227 725
rect 5130 634 5136 719
rect 5136 634 5221 719
rect 5221 634 5227 719
rect 5130 628 5227 634
rect 5440 592 5537 760
rect 5927 568 6016 760
rect 6924 636 7032 642
rect 6924 540 6930 636
rect 6930 540 7026 636
rect 7026 540 7032 636
rect 6924 534 7032 540
rect 7272 492 7380 684
rect 172 182 224 246
rect 5326 189 5378 241
rect 1991 -133 2065 -81
<< metal2 >>
rect 296 10920 382 10926
rect -53 10793 -47 10879
rect 39 10793 296 10879
rect 296 10746 382 10752
rect 130 10284 222 10290
rect 306 10200 312 10322
rect 480 10200 486 10322
rect 130 9252 222 10192
rect 335 9913 457 10200
rect 335 9791 4375 9913
rect 2376 9326 2536 9332
rect 130 9162 2250 9252
rect 130 9160 2256 9162
rect 2152 9040 2256 9160
rect 2367 9134 2376 9326
rect 2376 9128 2536 9134
rect 160 9000 224 9006
rect 2114 9000 2120 9040
rect 224 8936 2120 9000
rect 160 8930 224 8936
rect 2114 8872 2120 8936
rect 2288 9000 2294 9040
rect 2288 8936 4042 9000
rect 2288 8872 2294 8936
rect 672 8824 864 8833
rect 666 8766 672 8824
rect 864 8766 870 8824
rect 672 8759 864 8766
rect 306 8488 396 8494
rect -5 8359 1 8449
rect 91 8359 306 8449
rect 1986 8320 1992 8384
rect 2056 8320 2062 8384
rect 306 8314 396 8320
rect 1995 8138 2054 8320
rect 1960 8046 1982 8138
rect 2074 8046 2088 8138
rect 3978 3970 4042 8936
rect 4253 8301 4375 9791
rect 4253 8173 4375 8179
rect 3978 3900 4042 3906
rect 5440 3162 5552 3168
rect 5088 3022 5094 3134
rect 5206 3022 5440 3134
rect 5440 2988 5552 2994
rect 5308 2532 5372 2538
rect 5308 2172 5372 2468
rect 6108 2172 6172 2178
rect 5308 2108 6108 2172
rect 6108 2102 6172 2108
rect 5440 2014 5535 2020
rect 5099 1871 5105 1966
rect 5200 1871 5440 1966
rect 5440 1816 5535 1822
rect 7272 1826 7350 1832
rect 6975 1703 6981 1781
rect 7059 1703 7272 1781
rect 7272 1652 7350 1658
rect 288 760 389 766
rect -36 626 -30 727
rect 71 626 288 727
rect 5440 760 5537 766
rect 288 586 389 592
rect 2695 630 2747 636
rect 5124 628 5130 725
rect 5227 628 5440 725
rect 5440 586 5537 592
rect 5927 760 6016 766
rect 2695 572 2747 578
rect 172 246 224 252
rect 2698 237 2743 572
rect 6016 620 6634 709
rect 7272 684 7380 690
rect 6945 642 7034 650
rect 5927 562 6016 568
rect 6545 605 6634 620
rect 6918 605 6924 642
rect 6545 534 6924 605
rect 7032 534 7272 642
rect 6545 516 7034 534
rect 7272 486 7380 492
rect 5320 237 5326 241
rect 224 192 5326 237
rect 1987 190 2032 192
rect 5320 189 5326 192
rect 5378 189 5384 241
rect 172 176 224 182
rect 1982 -133 1991 -59
rect 2065 -133 2074 -59
rect 1991 -139 2065 -133
<< via2 >>
rect 2376 9134 2498 9326
rect 672 8768 864 8824
rect 1982 8046 2074 8138
rect 1991 -81 2065 -59
rect 1991 -133 2065 -81
<< metal3 >>
rect 2371 9326 2503 9331
rect 2371 9296 2376 9326
rect 630 9164 2376 9296
rect 2371 9134 2376 9164
rect 2498 9134 2503 9326
rect 2371 9129 2503 9134
rect 667 8829 869 8835
rect 667 8759 869 8765
rect 1977 8138 2079 8143
rect 1977 8046 1982 8138
rect 2074 8046 2079 8138
rect 1977 8041 2079 8046
rect 1986 -59 2070 8041
rect 1986 -133 1991 -59
rect 2065 -133 2070 -59
rect 1986 -138 2070 -133
<< via3 >>
rect 667 8824 869 8829
rect 667 8768 672 8824
rect 672 8768 864 8824
rect 864 8768 869 8824
rect 667 8765 869 8768
<< metal4 >>
rect 738 8830 798 9140
rect 666 8829 870 8830
rect 666 8765 667 8829
rect 869 8765 870 8829
rect 666 8764 870 8765
use JNWATR_PCH_4C1F2  xa1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWTR_RPPO16  xa2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1743091282
transform 1 0 0 0 1 978
box 0 0 4472 3440
use JNWTR_RPPO16  xa3
timestamp 1743091282
transform 1 0 0 0 1 4682
box 0 0 4472 3440
use JNWATR_PCH_4C1F2  xb1
timestamp 1734044400
transform 1 0 5152 0 1 0
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xb2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5152 0 1 1326
box -184 -128 1336 928
use JNWATR_NCH_4C1F2  xb3 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5152 0 1 2402
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xc2
timestamp 1734044400
transform 1 0 6984 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C1F2  xc3
timestamp 1734044400
transform 1 0 6984 0 1 1066
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xd
timestamp 1734044400
transform 1 0 0 0 1 8280
box -184 -128 1336 928
use JNWTR_CAPX1  xd1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1723932000
transform 1 0 0 0 1 9080
box 0 0 1080 1080
use JNWATR_NCH_4C1F2  xd2
timestamp 1734044400
transform 1 0 0 0 1 10160
box -184 -128 1336 928
use JNWATR_NCH_2C1F2  xe ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 1832 0 1 8280
box -184 -128 1208 928
<< labels >>
flabel metal1 5404 6258 5806 6676 0 FreeSans 800 0 0 0 VSS
flabel metal1 2664 -72 3074 130 0 FreeSans 800 0 0 0 VDD
flabel metal1 4740 1048 4922 1206 0 FreeSans 800 0 0 0 VIN-
flabel metal1 6594 30 6764 220 0 FreeSans 800 0 0 0 VIN+
flabel metal1 1450 9330 1756 9598 0 FreeSans 800 0 0 0 VOUT
<< properties >>
string FIXED_BBOX 0 0 8136 10960
<< end >>
