magic
tech sky130A
magscale 1 2
timestamp 1744208368
<< error_s >>
rect 16415 12249 16652 12269
rect 16435 12230 16436 12249
rect 16632 12230 16652 12249
<< viali >>
rect 15704 11180 15884 11372
rect 364 5906 604 6078
rect 3912 5906 4108 6146
rect 4356 3012 4456 3124
rect 484 2474 584 2574
rect 3870 2438 4042 2610
rect 4344 -464 4456 -364
<< metal1 >>
rect 3657 14069 3928 14075
rect 3657 13868 3928 13874
rect 18113 12118 18552 12198
rect 15960 12054 18552 12118
rect 15960 11904 16024 12054
rect 15754 11876 15882 11882
rect 15754 11742 15882 11748
rect 16082 11716 16088 11908
rect 16216 11716 16222 11908
rect 16472 11844 16664 11850
rect 18113 11813 18552 12054
rect 18206 11812 18552 11813
rect 16472 11714 16664 11720
rect 15698 11378 15890 11384
rect 15692 11174 15698 11378
rect 15867 11372 15890 11378
rect 15884 11180 15890 11372
rect 16491 11301 17218 11456
rect 17373 11301 17379 11456
rect 15867 11174 15890 11180
rect 15698 11168 15890 11174
rect 4726 6650 4949 6656
rect 1608 6427 4726 6650
rect 4726 6421 4949 6427
rect 21213 6460 21677 6466
rect 21213 6237 21677 6243
rect 3906 6146 4114 6158
rect 352 6078 616 6084
rect 352 5906 364 6078
rect 604 5906 616 6078
rect 352 5900 616 5906
rect 3906 5906 3912 6146
rect 4108 6130 4114 6146
rect 5316 6136 5530 6142
rect 4108 5989 5316 6130
rect 5530 6130 5652 6136
rect 5530 5989 7814 6130
rect 4108 5922 7814 5989
rect 4108 5906 4114 5922
rect 392 4428 576 5900
rect 3906 5894 4114 5906
rect 392 4244 4048 4428
rect 3864 4010 4048 4244
rect 3858 3826 4054 4010
rect 3864 3533 4048 3826
rect 4189 3533 4323 3539
rect 3864 3399 4189 3533
rect 3864 2610 4048 3399
rect 4189 3393 4323 3399
rect 4350 3124 4462 3136
rect 4350 3012 4356 3124
rect 4456 3012 5540 3124
rect 4350 3000 4462 3012
rect 478 2574 590 2586
rect 478 2474 484 2574
rect 584 2474 590 2574
rect 478 650 590 2474
rect 3864 2438 3870 2610
rect 4042 2438 4048 2610
rect 3864 2426 4048 2438
rect 5428 650 5540 3012
rect 7606 2033 7814 5922
rect 10344 4715 10350 4934
rect 10569 4715 10575 4934
rect 10350 4094 10569 4715
rect 10816 4194 10822 4418
rect 11046 4194 11052 4418
rect 10822 4094 11046 4194
rect 10350 3875 11046 4094
rect 10822 2048 11046 3875
rect 7359 1533 7907 2033
rect 10146 1798 11106 2048
rect 478 538 5540 650
rect 5428 -358 5540 538
rect 7472 -4 7640 1533
rect 10128 1318 11106 1798
rect 7466 -172 7472 -4
rect 7640 -172 7646 -4
rect 10532 -358 10644 1318
rect 20526 1038 20532 1228
rect 20682 1038 20688 1228
rect 22388 1069 22394 1224
rect 22549 1069 22555 1224
rect 22394 246 22549 1069
rect 22383 240 22549 246
rect 22394 68 22549 240
rect 22383 62 22549 68
rect 22394 59 22549 62
rect 16344 -172 16350 -4
rect 16518 -172 16524 -4
rect 4332 -364 10644 -358
rect 4332 -464 4344 -364
rect 4456 -464 10644 -364
rect 4332 -470 10644 -464
<< via1 >>
rect 3657 13874 3928 14069
rect 15754 11748 15882 11876
rect 16088 11716 16216 11908
rect 16472 11720 16664 11844
rect 15698 11372 15867 11378
rect 15698 11180 15704 11372
rect 15704 11180 15867 11372
rect 17218 11301 17373 11456
rect 15698 11174 15867 11180
rect 4726 6427 4949 6650
rect 21213 6243 21677 6460
rect 5316 5989 5530 6136
rect 4189 3399 4323 3533
rect 10350 4715 10569 4934
rect 10822 4194 11046 4418
rect 7472 -172 7640 -4
rect 20532 1038 20682 1228
rect 22394 1069 22549 1224
rect 16350 -172 16518 -4
<< metal2 >>
rect 875 16075 16632 16272
rect 875 15887 1072 16075
rect 3651 13874 3657 14069
rect 3928 13874 3934 14069
rect 3657 13865 3928 13874
rect 16435 12249 16632 16075
rect 16435 12052 16632 12062
rect 16088 11908 16216 11914
rect 15748 11748 15754 11876
rect 15882 11748 16088 11876
rect 16472 11844 16664 11853
rect 16466 11720 16472 11844
rect 16664 11720 16670 11844
rect 16088 11710 16216 11716
rect 17218 11456 17373 11462
rect 15698 11378 15867 11384
rect 15689 11174 15698 11378
rect 17373 11301 17382 11456
rect 17218 11295 17373 11301
rect 15698 11168 15867 11174
rect 4720 6427 4726 6650
rect 4949 6427 4955 6650
rect 21213 6460 21677 6466
rect 4728 4934 4947 6427
rect 21207 6243 21213 6460
rect 21677 6243 21683 6460
rect 21213 6234 21677 6243
rect 5316 6136 5530 6145
rect 5310 5989 5316 6136
rect 5530 5989 5536 6136
rect 10350 4934 10569 4940
rect 4728 4715 10350 4934
rect 10822 4809 11046 4814
rect 10350 4709 10569 4715
rect 10818 4595 10827 4809
rect 11041 4595 11050 4809
rect 10822 4418 11046 4595
rect 10822 4188 11046 4194
rect 4644 3533 4768 3537
rect 4183 3399 4189 3533
rect 4323 3528 4773 3533
rect 4323 3404 4644 3528
rect 4768 3404 4773 3528
rect 4323 3399 4773 3404
rect 4644 3395 4768 3399
rect 22394 1509 22549 1514
rect 22390 1364 22399 1509
rect 22544 1364 22553 1509
rect 20532 1228 20682 1234
rect 20523 1038 20532 1228
rect 22394 1224 22549 1364
rect 22394 1063 22549 1069
rect 20532 1032 20682 1038
rect 7472 -4 7640 2
rect 16350 -4 16518 2
rect 7640 -172 16350 -4
rect 7472 -178 7640 -172
rect 16350 -178 16518 -172
<< via2 >>
rect 3657 13874 3928 14059
rect 16435 12062 16632 12249
rect 16472 11730 16664 11844
rect 15698 11174 15843 11378
rect 17228 11301 17373 11456
rect 21213 6243 21677 6457
rect 5316 6021 5530 6136
rect 10827 4595 11041 4809
rect 4644 3404 4768 3528
rect 22399 1364 22544 1509
rect 20532 1038 20663 1228
<< metal3 >>
rect 3652 14062 3933 14068
rect 3652 13863 3933 13869
rect 16506 12254 16630 12380
rect 16430 12249 16637 12254
rect 16430 12062 16435 12249
rect 16632 12062 16637 12249
rect 16430 12057 16637 12062
rect 16506 11849 16630 12057
rect 16467 11844 16669 11849
rect 16467 11730 16472 11844
rect 16664 11730 16669 11844
rect 16467 11725 16669 11730
rect 15687 11169 15693 11383
rect 15846 11169 15852 11383
rect 17219 11296 17225 11461
rect 17378 11296 17384 11461
rect 21208 6460 21682 6466
rect 21208 6232 21682 6238
rect 5311 6141 5535 6147
rect 5311 6021 5316 6037
rect 5530 6021 5535 6037
rect 5311 6016 5535 6021
rect 10822 5171 11046 5172
rect 10817 4949 10823 5171
rect 11045 4949 11051 5171
rect 10822 4809 11046 4949
rect 10822 4595 10827 4809
rect 11041 4595 11046 4809
rect 10822 4590 11046 4595
rect 4926 3533 5058 3538
rect 4639 3532 5059 3533
rect 4639 3528 4926 3532
rect 4639 3404 4644 3528
rect 4768 3404 4926 3528
rect 4639 3400 4926 3404
rect 5058 3400 5059 3532
rect 4639 3399 5059 3400
rect 4926 3394 5058 3399
rect 22394 1935 22549 1936
rect 22389 1782 22395 1935
rect 22548 1782 22554 1935
rect 22394 1509 22549 1782
rect 22394 1364 22399 1509
rect 22544 1364 22549 1509
rect 22394 1359 22549 1364
rect 20521 1033 20527 1233
rect 20659 1228 20668 1233
rect 20663 1038 20668 1228
rect 20659 1033 20668 1038
<< via3 >>
rect 3652 14059 3933 14062
rect 3652 13874 3657 14059
rect 3657 13874 3928 14059
rect 3928 13874 3933 14059
rect 3652 13869 3933 13874
rect 15693 11378 15846 11383
rect 15693 11174 15698 11378
rect 15698 11174 15843 11378
rect 15843 11174 15846 11378
rect 15693 11169 15846 11174
rect 17225 11456 17378 11461
rect 17225 11301 17228 11456
rect 17228 11301 17373 11456
rect 17373 11301 17378 11456
rect 17225 11296 17378 11301
rect 21208 6457 21682 6460
rect 21208 6243 21213 6457
rect 21213 6243 21677 6457
rect 21677 6243 21682 6457
rect 21208 6238 21682 6243
rect 5311 6136 5535 6141
rect 5311 6037 5316 6136
rect 5316 6037 5530 6136
rect 5530 6037 5535 6136
rect 10823 4949 11045 5171
rect 4926 3400 5058 3532
rect 22395 1782 22548 1935
rect 20527 1228 20659 1233
rect 20527 1038 20532 1228
rect 20532 1038 20659 1228
rect 20527 1033 20659 1038
<< metal4 >>
rect 3651 14062 3934 14063
rect 3651 13869 3652 14062
rect 3933 13869 3934 14062
rect 3651 13868 3934 13869
rect 3695 6962 3890 13868
rect 15496 12190 15888 12250
rect 15496 11354 15556 12190
rect 17224 11461 17379 11462
rect 15692 11383 15847 11384
rect 15692 11354 15693 11383
rect 15427 11199 15693 11354
rect 3695 6767 5510 6962
rect 5354 6142 5492 6767
rect 5310 6141 5536 6142
rect 5310 6037 5311 6141
rect 5535 6037 5536 6141
rect 5310 6036 5536 6037
rect 5354 6020 5492 6036
rect 15427 5172 15582 11199
rect 15692 11169 15693 11199
rect 15846 11169 15847 11383
rect 17224 11296 17225 11461
rect 17378 11456 17379 11461
rect 17378 11301 22549 11456
rect 17378 11296 17379 11301
rect 17224 11295 17379 11296
rect 15692 11168 15847 11169
rect 21207 6460 21683 6461
rect 21207 6238 21208 6460
rect 21682 6238 21683 6460
rect 21207 6237 21683 6238
rect 21333 5172 21557 6237
rect 10822 5171 21557 5172
rect 10822 4949 10823 5171
rect 11045 4949 21557 5171
rect 10822 4948 21557 4949
rect 4925 3532 5059 3533
rect 4925 3400 4926 3532
rect 5058 3400 5059 3532
rect 4925 1200 5059 3400
rect 22394 1935 22549 11301
rect 22394 1782 22395 1935
rect 22548 1782 22549 1935
rect 22394 1781 22549 1782
rect 20526 1233 20660 1234
rect 20526 1200 20527 1233
rect 4925 1066 20527 1200
rect 20526 1033 20527 1066
rect 20659 1033 20660 1233
rect 20526 1032 20660 1033
use JNWTR_RPPO16  xa2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1743091282
transform 1 0 0 0 1 -512
box 0 0 4472 3440
use JNWTR_RPPO16  xa3
timestamp 1743091282
transform 1 0 0 0 1 2986
box 0 0 4472 3440
use temo_effected_current  xa4 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_GR01_SKY130A
timestamp 1744202613
transform 1 0 0 0 1 6880
box -184 -472 15120 9410
use SKYOP  xb1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_GR01_SKY130A
timestamp 1744207573
transform 1 0 15800 0 1 0
box -184 -178 8320 11088
use JNWATR_NCH_4C5F0  xb2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 15800 0 1 11220
box -184 -128 1336 928
use JNWTR_CAPX1  xb3 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1723932000
transform 1 0 15800 0 1 12190
box 0 0 1080 1080
<< labels >>
flabel metal1 7384 1558 7870 2010 0 FreeSans 800 0 0 0 VDD
flabel metal1 10172 1352 11062 1956 0 FreeSans 800 0 0 0 VSS
flabel metal1 18140 11834 18526 12170 0 FreeSans 800 0 0 0 reset
flabel space 17262 9332 17586 9598 0 FreeSans 1600 0 0 0 cmp
<< properties >>
string FIXED_BBOX 0 0 23936 15800
<< end >>
