*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/aop_v4_lpe.spi
#else
.include ../../../work/xsch/aop_v4.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS   dc  {AVDD}


VIN+ IN+ VIN_OFFSET+ dc 0 sin (0 10m 1Meg 0 0 0)
VIN- IN- VIN_OFFSET- dc 0 sin (0 10m 1Meg 0 0 180)
VOFFP VIN_OFFSET+ VSS dc  0.81
V0FFp VIN_OFFSET- VSS dc 0.81
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.save @r.xdut.R1[i]

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit
optran 0 0 0 1n 1u 0

*dc temp -60 120 1
tran 1n 10u 1p
write
quit


.endc

.end
