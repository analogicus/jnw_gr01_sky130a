magic
tech sky130A
magscale 1 2
timestamp 1744390707
<< locali >>
rect 10440 3624 11604 3640
rect 10552 3528 11604 3624
<< viali >>
rect -95 9687 68 9850
rect 9298 6463 9499 6664
rect 11028 6463 11268 6672
rect 10440 3528 10552 3624
rect 9302 2966 9482 3146
rect 9764 2959 10004 3160
rect 6992 2212 7232 2440
rect 9178 -8 9317 131
rect 10228 26 10324 122
<< metal1 >>
rect 1926 11784 2828 11950
rect 672 11592 2828 11784
rect 160 11028 224 11344
rect 288 10800 480 11464
rect 1918 11378 2828 11592
rect 4374 11280 5146 11281
rect 160 10228 224 10508
rect 288 10056 480 10746
rect 4074 10724 5346 11280
rect 676 10503 6121 10724
rect 4074 10490 5346 10503
rect -101 9856 74 9862
rect -101 9675 74 9681
rect 299 9672 305 9864
rect 480 9672 486 9864
rect 160 8266 224 9672
rect 688 9198 841 9778
rect 688 9039 841 9045
rect 160 8202 2750 8266
rect 5900 7340 6121 10503
rect 5900 7119 11259 7340
rect 5502 6819 5508 6846
rect 4693 6677 4699 6819
rect 4841 6677 5508 6819
rect 5502 6671 5508 6677
rect 5683 6819 5689 6846
rect 6596 6819 7584 6962
rect 5683 6677 7584 6819
rect 11038 6678 11259 7119
rect 5683 6671 5689 6677
rect 6596 6438 7584 6677
rect 9292 6664 9505 6676
rect 9292 6463 9298 6664
rect 9499 6463 9505 6664
rect 6596 6436 6749 6438
rect 3021 3601 3233 3719
rect 3351 3601 3357 3719
rect 3021 2717 3139 3601
rect 6992 2446 7232 6438
rect 9292 5452 9505 6463
rect 11016 6672 11280 6678
rect 11016 6463 11028 6672
rect 11268 6463 11280 6672
rect 11016 6457 11280 6463
rect 9292 5239 9991 5452
rect 9778 3547 9991 5239
rect 10428 3624 10564 3630
rect 9772 3328 9778 3547
rect 9991 3328 9997 3547
rect 10428 3528 10440 3624
rect 10552 3528 10564 3624
rect 10428 3522 10564 3528
rect 9778 3166 9991 3328
rect 9752 3160 10016 3166
rect 7376 3146 9494 3152
rect 7376 2966 9302 3146
rect 9482 2966 9494 3146
rect 7376 2960 9494 2966
rect 6980 2440 7244 2446
rect 6980 2212 6992 2440
rect 7232 2212 7244 2440
rect 6980 2206 7244 2212
rect 7376 1776 7568 2960
rect 9752 2959 9764 3160
rect 10004 2959 10016 3160
rect 9752 2953 10016 2959
rect 7248 1160 7312 1392
rect 7760 976 7952 1556
rect 4777 797 4783 959
rect 4945 797 4951 959
rect 4783 541 4945 797
rect 7370 662 7376 854
rect 7529 662 7535 854
rect 7248 28 7312 584
rect 4898 4 7312 28
rect 7760 4 7952 750
rect 9172 131 9323 143
rect 4898 -135 8332 4
rect 9172 -8 9178 131
rect 9317 -8 9323 131
rect 10442 128 10550 3522
rect 10216 122 10550 128
rect 10216 26 10228 122
rect 10324 26 10550 122
rect 10216 20 10550 26
rect 9172 -135 9323 -8
rect 4898 -212 9323 -135
rect 6723 -286 9323 -212
rect 6723 -426 8332 -286
<< via1 >>
rect -101 9850 74 9856
rect -101 9687 -95 9850
rect -95 9687 68 9850
rect 68 9687 74 9850
rect -101 9681 74 9687
rect 305 9672 480 9864
rect 688 9045 841 9198
rect 4699 6677 4841 6819
rect 5508 6671 5683 6846
rect 3233 3601 3351 3719
rect 9778 3328 9991 3547
rect 4783 797 4945 959
rect 7376 662 7529 854
<< metal2 >>
rect 305 9864 480 9870
rect -107 9681 -101 9856
rect 74 9681 305 9856
rect 480 9681 5683 9856
rect 305 9666 480 9672
rect 682 9045 688 9198
rect 841 9045 5129 9198
rect 4699 6819 4841 7049
rect 4699 6671 4841 6677
rect 4976 5418 5129 9045
rect 5508 6846 5683 9681
rect 5508 6665 5683 6671
rect 4976 5265 6811 5418
rect 3221 3931 3364 3940
rect 6658 3939 6811 5265
rect 3221 3779 3364 3788
rect 6649 3780 6658 3939
rect 6801 3780 6811 3939
rect 3233 3719 3351 3779
rect 3233 3595 3351 3601
rect 4783 3488 4945 3493
rect 4755 3336 4764 3488
rect 4965 3336 4974 3488
rect 4783 959 4945 3336
rect 4783 791 4945 797
rect 6658 835 6811 3780
rect 9778 3547 9991 3553
rect 9769 3328 9778 3547
rect 9778 3322 9991 3328
rect 7376 854 7529 860
rect 6658 682 7376 835
rect 7376 656 7529 662
<< via2 >>
rect 3221 3788 3364 3931
rect 6658 3780 6801 3939
rect 4764 3336 4965 3488
rect 9778 3328 9981 3547
<< metal3 >>
rect 6653 3939 6806 3944
rect 6653 3936 6658 3939
rect 3216 3931 6658 3936
rect 3216 3788 3221 3931
rect 3364 3788 6658 3931
rect 3216 3783 6658 3788
rect 6653 3780 6658 3783
rect 6801 3780 6806 3939
rect 6653 3775 6806 3780
rect 4759 3492 4970 3493
rect 4753 3332 4759 3492
rect 4970 3332 4976 3492
rect 4759 3331 4970 3332
rect 9767 3323 9773 3552
rect 9984 3323 9990 3552
<< via3 >>
rect 4759 3488 4970 3492
rect 4759 3336 4764 3488
rect 4764 3336 4965 3488
rect 4965 3336 4970 3488
rect 4759 3332 4970 3336
rect 9773 3547 9984 3552
rect 9773 3328 9778 3547
rect 9778 3328 9981 3547
rect 9981 3328 9984 3547
rect 9773 3323 9984 3328
<< metal4 >>
rect 9772 3552 9985 3553
rect 9772 3544 9773 3552
rect 4758 3492 9773 3544
rect 4758 3332 4759 3492
rect 4970 3332 9773 3492
rect 4758 3331 9773 3332
rect 9772 3323 9773 3331
rect 9984 3323 9985 3552
rect 9772 3322 9985 3323
use SKY_OTA  xa2
timestamp 1744388539
transform 1 0 0 0 1 0
box -184 -460 6592 8906
use JNWATR_PCH_4C5F0  xb1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 7088 0 1 480
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xb2
timestamp 1740610800
transform 1 0 7088 0 1 1280
box -184 -128 1336 928
use JNWTR_RPPO2  xc1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744368746
transform 1 0 8920 0 1 0
box 0 0 1448 3440
use JNWTR_RPPO8  xc2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744286843
transform 1 0 8920 0 1 3512
box 0 0 2744 3440
use JNWATR_PCH_4C5F0  xe1
timestamp 1740610800
transform 1 0 0 0 1 9560
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xe2
timestamp 1740610800
transform 1 0 0 0 1 10360
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xe3
timestamp 1740610800
transform 1 0 0 0 1 11160
box -184 -128 1336 928
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT0 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 7088 0 1 0
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT2
timestamp 1740610800
transform 1 0 0 0 1 9080
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 7088 0 1 2080
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP3
timestamp 1740610800
transform 1 0 0 0 1 11960
box -184 -128 1336 608
<< labels >>
flabel metal1 6660 6480 7534 6902 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 6804 -362 8306 -42 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 4128 10534 5270 11202 0 FreeSans 1600 0 0 0 Vref
port 3 nsew
flabel metal1 1978 11428 2782 11892 0 FreeSans 1600 0 0 0 OUT
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 11664 12440
<< end >>
