magic
tech sky130A
magscale 1 2
timestamp 1744202613
<< viali >>
rect 1780 8828 1905 8953
rect -67 8661 36 8764
rect 3616 8650 3741 8775
rect 11045 6477 11243 6675
rect 14516 6464 14756 6692
rect 14992 3548 15104 3648
rect 14998 3266 15098 3366
rect 11016 2926 11196 3106
rect 14516 2962 14756 3160
rect 8720 1464 8912 1616
rect 11100 -66 11280 114
<< metal1 >>
rect 160 9398 2052 9410
rect 160 9346 3886 9398
rect 160 8816 224 9346
rect 1988 9334 3886 9346
rect 1988 8978 2052 9334
rect 1774 8959 1911 8965
rect 672 8846 864 8852
rect -73 8770 42 8776
rect -73 8649 42 8655
rect 282 8616 288 8808
rect 403 8616 409 8808
rect 1774 8816 1911 8822
rect 2114 8794 2120 8986
rect 2257 8794 2263 8986
rect 3822 8808 3886 9334
rect 672 8761 864 8767
rect 3610 8781 3747 8787
rect 3610 8638 3747 8644
rect 3946 8616 3952 8808
rect 4089 8616 4095 8808
rect 160 6852 224 8224
rect 324 8002 444 8388
rect 2120 8002 2312 8614
rect 2504 8516 2696 8522
rect 2504 8348 2696 8354
rect 324 7882 2312 8002
rect 3952 7886 4144 8424
rect 2120 7844 2312 7882
rect 3694 7694 4144 7886
rect 4310 7242 4550 8370
rect 4310 7002 14756 7242
rect 160 6788 830 6852
rect 14516 6698 14756 7002
rect 14504 6692 14768 6698
rect 11039 6675 11249 6687
rect 11039 6477 11045 6675
rect 11243 6477 11249 6675
rect 11039 5201 11249 6477
rect 14504 6464 14516 6692
rect 14756 6464 14768 6692
rect 14504 6458 14768 6464
rect 11039 4991 14741 5201
rect 14531 3557 14741 4991
rect 14980 3648 15116 3654
rect 14525 3347 14531 3557
rect 14741 3347 14747 3557
rect 14980 3548 14992 3648
rect 15104 3548 15116 3648
rect 14980 3542 15116 3548
rect 14992 3366 15104 3542
rect 14531 3166 14741 3347
rect 14992 3266 14998 3366
rect 15098 3266 15104 3366
rect 14992 3254 15104 3266
rect 14504 3160 14768 3166
rect 9104 3106 11208 3112
rect 9104 2926 11016 3106
rect 11196 2926 11208 3106
rect 14504 2962 14516 3160
rect 14756 2962 14768 3160
rect 14504 2956 14768 2962
rect 9104 2920 11208 2926
rect 7280 2254 7444 2260
rect 7280 2084 7444 2090
rect 8714 1622 8918 1628
rect 8708 1458 8714 1622
rect 8918 1458 8924 1622
rect 8714 1452 8918 1458
rect 9104 1200 9296 2920
rect 4711 1158 4858 1164
rect 4711 1005 4858 1011
rect 8976 660 9040 916
rect 9488 542 9680 1072
rect 9145 404 9277 410
rect 9145 251 9277 257
rect 7727 -205 7854 -199
rect 6934 -382 6998 -244
rect 7445 -332 7727 -205
rect 7727 -338 7854 -332
rect 8976 -280 9040 108
rect 9488 -280 9680 232
rect 11094 114 11286 126
rect 11094 -66 11100 114
rect 11280 -66 11286 114
rect 11094 -280 11286 -66
rect 8976 -382 11286 -280
rect 6934 -446 11286 -382
rect 8976 -472 11286 -446
<< via1 >>
rect 1774 8953 1911 8959
rect -73 8764 42 8770
rect -73 8661 -67 8764
rect -67 8661 36 8764
rect 36 8661 42 8764
rect -73 8655 42 8661
rect 288 8616 403 8808
rect 672 8767 864 8846
rect 1774 8828 1780 8953
rect 1780 8828 1905 8953
rect 1905 8828 1911 8953
rect 1774 8822 1911 8828
rect 2120 8794 2257 8986
rect 3610 8775 3747 8781
rect 3610 8650 3616 8775
rect 3616 8650 3741 8775
rect 3741 8650 3747 8775
rect 3610 8644 3747 8650
rect 3952 8616 4089 8808
rect 2504 8354 2696 8516
rect 14531 3347 14741 3557
rect 7280 2090 7444 2254
rect 8714 1616 8918 1622
rect 8714 1464 8720 1616
rect 8720 1464 8912 1616
rect 8912 1464 8918 1616
rect 8714 1458 8918 1464
rect 4711 1011 4858 1158
rect 9145 257 9277 404
rect 7727 -332 7854 -205
<< metal2 >>
rect 729 9120 1103 9235
rect 732 9065 1103 9120
rect 729 8975 1103 9065
rect 2120 8986 2257 8992
rect 729 8846 808 8975
rect 288 8808 403 8814
rect -79 8655 -73 8770
rect 42 8655 288 8770
rect 666 8767 672 8846
rect 864 8767 870 8846
rect 1768 8822 1774 8959
rect 1911 8822 2120 8959
rect 2120 8788 2257 8794
rect 3952 8808 4089 8814
rect 3604 8644 3610 8781
rect 3747 8644 3952 8781
rect 288 8610 403 8616
rect 3952 8610 4089 8616
rect 2498 8354 2504 8516
rect 2696 8354 2702 8516
rect 2504 8345 2696 8354
rect 14531 3557 14741 3563
rect 10287 3347 14531 3557
rect 7274 2090 7280 2254
rect 7444 2090 8898 2254
rect 8734 1622 8898 2090
rect 8708 1458 8714 1622
rect 8918 1458 8924 1622
rect 4711 1158 4858 1167
rect 4705 1011 4711 1158
rect 4858 1011 4864 1158
rect 4711 1002 4858 1011
rect 9130 404 9277 413
rect 9277 257 9283 404
rect 9130 248 9277 257
rect 10320 -205 10465 3347
rect 14531 3341 14741 3347
rect 7721 -332 7727 -205
rect 7854 -332 10465 -205
rect 10320 -342 10465 -332
<< via2 >>
rect 2504 8354 2696 8501
rect 4711 1011 4858 1158
rect 9130 257 9145 404
rect 9145 257 9277 404
<< metal3 >>
rect 2499 8501 2701 8506
rect 2499 8354 2504 8501
rect 2696 8354 2701 8501
rect 2499 8349 2701 8354
rect 2522 7961 2679 8349
rect 2522 7804 4954 7961
rect 4797 5075 4954 7804
rect 4797 4918 8544 5075
rect 8387 1163 8544 4918
rect 4706 1158 8544 1163
rect 4706 1011 4711 1158
rect 4858 1011 8544 1158
rect 4706 1006 8544 1011
rect 8387 409 8544 1006
rect 8387 404 9282 409
rect 8387 257 9130 404
rect 9277 257 9282 404
rect 8387 252 9282 257
use SKY_OTA  xa2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_GR01_SKY130A
timestamp 1744189113
transform 1 0 0 0 1 0
box -184 -453 8320 7964
use JNWATR_PCH_4C5F0  xb1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 8816 0 1 0
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xb2
timestamp 1734044400
transform 1 0 8816 0 1 800
box -184 -128 1336 928
use JNWTR_RPPO16  xc1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1743091282
transform 1 0 10648 0 1 0
box 0 0 4472 3440
use JNWTR_RPPO16  xc2
timestamp 1743091282
transform 1 0 10648 0 1 3532
box 0 0 4472 3440
use JNWATR_PCH_4C5F0  xd1
timestamp 1734044400
transform 1 0 0 0 1 8120
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xe1
timestamp 1734044400
transform 1 0 1832 0 1 8310
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xf
timestamp 1734044400
transform 1 0 3664 0 1 8120
box -184 -128 1336 928
<< labels >>
flabel space 3686 7030 3892 7282 0 FreeSans 800 0 0 0 VDD
flabel space 1622 -438 1828 -186 0 FreeSans 800 0 0 0 VSS
flabel metal2 744 8982 1084 9214 0 FreeSans 800 0 0 0 OUT
<< properties >>
string FIXED_BBOX 0 0 15120 8920
<< end >>
