*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/temo_effected_current_lpe.spi
#else
.include ../../../work/xsch/temo_effected_current.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
*.param TRF = 10p
*.param AVDD = {vdda}
.param TRF = 10p
.param AVDD = 1.8

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
*VSS  VSS  0     dc 0
*VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VSS  VSS  0     dc 0
VDD  VDD  0  dc {AVDD}
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.save all
.save i(v.xdut.v2)
.save v(xdut.vr) v(VDD) v(VSS) v(xdut.right_side)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit



optran 0 0 0 5n 80u 0

*dc temp -60 150 5
*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )


tran 1n 10n 1p
write
quit


.endc

.end
