magic
tech sky130A
magscale 1 2
timestamp 1744189113
<< locali >>
rect 1933 6834 1967 7309
rect 836 4338 896 4344
rect 836 4290 842 4338
rect 890 4290 896 4338
rect 836 4166 896 4290
rect 463 3942 604 3960
rect 467 3912 604 3942
rect 3949 3801 4027 3977
rect 467 3720 604 3732
rect 616 3440 2578 3496
rect 5329 1971 5371 2413
rect 5329 1932 5940 1971
rect 5329 1930 5371 1932
rect 5901 1874 5940 1932
rect 5901 1838 5940 1840
rect 6888 1688 7080 2302
rect 7139 1419 7202 1880
rect 5056 648 5248 1034
rect 5056 57 5248 152
rect 6922 60 7047 119
rect -93 -148 93 43
rect 5235 2 5248 57
rect -93 -183 -3 -148
rect 32 -183 93 -148
rect -93 -220 93 -183
rect 5056 -70 5248 2
rect -93 -275 95 -220
rect 5091 -158 5248 -70
rect 6888 -129 7080 60
rect 5091 -236 5252 -158
rect 6888 -184 6966 -129
rect 7021 -184 7080 -129
rect 6888 -194 7080 -184
rect 5091 -237 5300 -236
rect 5091 -262 5314 -237
rect -93 -341 93 -275
rect 5056 -304 5314 -262
rect 5056 -386 5300 -304
rect 5058 -404 5300 -386
rect 5233 -409 5300 -404
<< viali >>
rect 1664 7745 1856 7816
rect 1933 6800 1967 6834
rect 1664 5928 1856 6062
rect 842 4290 890 4338
rect 3949 3977 4027 4043
rect 428 3732 608 3912
rect 5056 2722 5248 2852
rect 6888 2302 7080 2482
rect 5830 1840 6010 1874
rect 7128 1880 7212 1964
rect 1374 844 1409 879
rect -3 -183 32 -148
rect 5056 -262 5091 -70
rect 6966 -184 7021 -129
rect 5314 -304 5369 -237
<< metal1 >>
rect 2048 7959 2240 7964
rect 1719 7899 2240 7959
rect 1719 7897 3767 7899
rect 1719 7876 3773 7897
rect 1719 7822 1802 7876
rect 2048 7837 3773 7876
rect 1652 7816 1868 7822
rect 1652 7745 1664 7816
rect 1856 7745 1868 7816
rect 1652 7739 1868 7745
rect 2048 7472 2240 7837
rect 738 6848 928 6888
rect 1905 6871 1991 6877
rect 1899 6865 1997 6871
rect 1146 6848 1206 6854
rect 738 6788 1146 6848
rect 738 6734 928 6788
rect 1146 6782 1206 6788
rect 1365 6770 1899 6865
rect 1365 6767 1997 6770
rect -164 6496 870 6560
rect 934 6496 940 6560
rect -164 4640 -100 6496
rect 1365 4781 1463 6767
rect 1899 6764 1997 6767
rect 1916 6560 1980 6566
rect 1916 6490 1980 6496
rect 2086 6454 2203 6764
rect 1652 6062 1868 6068
rect 1652 5928 1664 6062
rect 1856 5928 1868 6062
rect 1652 5922 1868 5928
rect 1690 5225 1831 5922
rect 2432 5885 2624 7304
rect 3691 7302 3773 7837
rect 3657 7087 3928 7302
rect 3656 6994 3928 7087
rect 3753 6755 3831 6994
rect 3753 6677 3949 6755
rect 4027 6677 4033 6755
rect 2432 5791 3041 5885
rect 3299 5791 3362 5797
rect 2432 5728 3299 5791
rect 2432 5699 3041 5728
rect 3299 5722 3362 5728
rect 2432 5696 2624 5699
rect 1690 5078 1831 5084
rect 2968 4987 3038 4993
rect 2968 4830 3038 4917
rect 1913 4828 4510 4830
rect 1913 4781 7848 4828
rect 1365 4683 7848 4781
rect -164 4576 224 4640
rect 1913 4636 7848 4683
rect 1913 4635 4510 4636
rect 160 534 224 4576
rect 830 4362 836 4422
rect 896 4362 902 4422
rect 5287 4377 5293 4507
rect 5423 4377 5429 4507
rect 836 4338 896 4362
rect 836 4290 842 4338
rect 890 4290 896 4338
rect 836 4278 896 4290
rect 3949 4361 4027 4367
rect 3949 4049 4027 4283
rect 3937 4043 4039 4049
rect 3937 3977 3949 4043
rect 4027 3977 4039 4043
rect 3937 3971 4039 3977
rect 416 3912 864 3918
rect 416 3732 428 3912
rect 608 3732 864 3912
rect 416 3726 864 3732
rect 672 175 864 3726
rect 5293 3362 5423 4377
rect 5093 3321 5632 3362
rect 5094 3306 5632 3321
rect 5094 3203 7080 3306
rect 5093 3170 7080 3203
rect 5093 2858 5211 3170
rect 5440 3114 7080 3170
rect 5044 2852 5260 2858
rect 5044 2722 5056 2852
rect 5248 2722 5260 2852
rect 5044 2716 5260 2722
rect 5440 2426 5632 3114
rect 6888 2734 7080 3114
rect 6888 2542 7464 2734
rect 6888 2488 7080 2542
rect 6876 2482 7092 2488
rect 6876 2302 6888 2482
rect 7080 2302 7092 2482
rect 6876 2296 7092 2302
rect 5824 1981 6016 2226
rect 5824 1970 6110 1981
rect 5824 1964 7224 1970
rect 5824 1880 7128 1964
rect 7212 1880 7224 1964
rect 5824 1874 7224 1880
rect 5824 1840 5830 1874
rect 6010 1864 6110 1874
rect 6010 1840 6016 1864
rect 5824 1506 6016 1840
rect 7272 1552 7464 2542
rect 7656 1540 7848 4636
rect 4692 1112 4884 1180
rect 4692 1048 5376 1112
rect 4692 1002 4884 1048
rect 4692 1000 4756 1002
rect 672 170 678 175
rect 156 111 229 117
rect 156 32 229 38
rect 666 -22 678 170
rect 749 111 864 175
rect 1368 879 1415 891
rect 1368 844 1374 879
rect 1409 844 1415 879
rect 749 38 838 111
rect 749 36 864 38
rect 749 -23 798 36
rect 1368 -142 1415 844
rect 5497 887 5583 1109
rect 5497 879 5963 887
rect 5497 801 7405 879
rect 5877 793 7405 801
rect 5877 611 5963 793
rect 7319 623 7405 793
rect 7656 568 7848 1274
rect 1468 38 1474 111
rect 1547 38 5378 111
rect 5050 -70 5097 -58
rect 1684 -142 1690 -89
rect -15 -148 1690 -142
rect -15 -183 -3 -148
rect 32 -183 1690 -148
rect -15 -189 1690 -183
rect 1555 -221 1690 -189
rect 1598 -230 1690 -221
rect 1831 -142 1837 -89
rect 5050 -142 5056 -70
rect 1831 -189 5056 -142
rect 1831 -230 1837 -189
rect 1598 -307 1831 -230
rect 5050 -262 5056 -189
rect 5091 -262 5097 -70
rect 7144 -60 7208 110
rect 6960 -129 7027 -117
rect 7144 -124 7542 -60
rect 6960 -184 6966 -129
rect 7021 -184 7027 -129
rect 5050 -274 5097 -262
rect 5308 -236 5375 -225
rect 6960 -236 7027 -184
rect 7478 -205 7542 -124
rect 5308 -237 7027 -236
rect 5308 -304 5314 -237
rect 5369 -303 7027 -237
rect 5369 -304 5375 -303
rect 1598 -340 1863 -307
rect 5308 -316 5375 -304
rect 7439 -333 7581 -205
rect 7463 -339 7581 -333
rect 1601 -353 1863 -340
rect 1601 -390 1864 -353
rect 1601 -453 1869 -390
<< via1 >>
rect 1146 6788 1206 6848
rect 1899 6834 1997 6865
rect 1899 6800 1933 6834
rect 1933 6800 1967 6834
rect 1967 6800 1997 6834
rect 1899 6770 1997 6800
rect 870 6496 934 6560
rect 1916 6496 1980 6560
rect 3949 6677 4027 6755
rect 3299 5728 3362 5791
rect 1690 5084 1831 5225
rect 2968 4917 3038 4987
rect 836 4362 896 4422
rect 5293 4377 5423 4507
rect 3949 4283 4027 4361
rect 156 38 229 111
rect 1474 38 1547 111
rect 1690 -230 1831 -89
<< metal2 >>
rect 1901 6870 1996 7413
rect 1330 6848 1386 6855
rect 1140 6788 1146 6848
rect 1206 6846 1388 6848
rect 1206 6790 1330 6846
rect 1386 6790 1388 6846
rect 1206 6788 1388 6790
rect 1330 6781 1386 6788
rect 1893 6770 1899 6865
rect 1997 6770 2003 6865
rect 3949 6755 4027 6761
rect 870 6560 934 6566
rect 934 6496 1916 6560
rect 1980 6496 1986 6560
rect 870 6490 934 6496
rect 3293 5728 3299 5791
rect 3362 5728 3368 5791
rect 3299 5532 3362 5728
rect 3293 5476 3302 5532
rect 3358 5476 3367 5532
rect 3299 5473 3362 5476
rect 1684 5084 1690 5225
rect 1831 5084 1837 5225
rect 836 4588 896 4590
rect 829 4532 838 4588
rect 894 4532 903 4588
rect 836 4422 896 4532
rect 836 4356 896 4362
rect 1474 111 1547 117
rect 150 38 156 111
rect 229 38 1474 111
rect 1474 32 1547 38
rect 1690 -89 1831 5084
rect 2968 4987 3038 4996
rect 2962 4917 2968 4987
rect 3038 4917 3044 4987
rect 3949 4475 4027 6677
rect 5293 4507 5423 4513
rect 3949 4409 5293 4475
rect 3949 4361 4027 4409
rect 5293 4371 5423 4377
rect 3943 4283 3949 4361
rect 4027 4283 4033 4361
rect 1690 -236 1831 -230
<< via2 >>
rect 1901 6865 1996 6870
rect 1330 6790 1386 6846
rect 1901 6785 1996 6865
rect 3302 5476 3358 5532
rect 838 4532 894 4588
rect 2968 4927 3038 4987
<< metal3 >>
rect 1901 6875 1996 7385
rect 1896 6870 2001 6875
rect 2065 6870 2160 6963
rect 1325 6846 1391 6851
rect 1325 6790 1330 6846
rect 1386 6790 1391 6846
rect 1325 6785 1391 6790
rect 1896 6785 1901 6870
rect 1996 6785 2321 6870
rect 1328 4900 1388 6785
rect 1896 6780 2321 6785
rect 1901 6775 2321 6780
rect 3297 5532 3363 5537
rect 3297 5476 3302 5532
rect 3358 5476 3363 5532
rect 3297 5471 3363 5476
rect 3298 5304 3361 5471
rect 3292 5251 3384 5304
rect 3271 5161 3277 5251
rect 3399 5161 3405 5251
rect 3292 5160 3384 5161
rect 2689 4987 3043 4992
rect 2689 4927 2968 4987
rect 3038 4927 3043 4987
rect 2689 4922 3043 4927
rect 1460 4902 1524 4908
rect 1002 4840 1460 4900
rect 1460 4832 1524 4838
rect 668 4592 732 4598
rect 833 4590 899 4593
rect 732 4588 899 4590
rect 732 4532 838 4588
rect 894 4532 899 4588
rect 732 4530 899 4532
rect 668 4522 732 4528
rect 833 4527 899 4530
<< via3 >>
rect 3277 5161 3399 5251
rect 1460 4838 1524 4902
rect 668 4528 732 4592
<< metal4 >>
rect 2776 5268 2841 5337
rect 3276 5251 3400 5252
rect 3276 5161 3277 5251
rect 3399 5161 3400 5251
rect 3276 4976 3400 5161
rect 1459 4902 1525 4903
rect 670 4593 730 4900
rect 1459 4838 1460 4902
rect 1524 4900 1525 4902
rect 1524 4840 1874 4900
rect 2782 4852 3400 4976
rect 1524 4838 1525 4840
rect 1459 4837 1525 4838
rect 667 4592 733 4593
rect 667 4528 668 4592
rect 732 4528 733 4592
rect 667 4527 733 4528
use JNWATR_NCH_4C5F0  xa1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 0 0 1 -130
box -184 -128 1336 928
use JNWTR_RPPO16  xa2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1743091282
transform 1 0 0 0 1 800
box 0 0 4472 3440
use JNWATR_NCH_4C5F0  xc1
timestamp 1734044400
transform 1 0 5152 0 1 0
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xc2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5152 0 1 2012
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xc3
timestamp 1734044400
transform 1 0 5152 0 1 938
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xd1
timestamp 1734044400
transform 1 0 6984 0 1 0
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xd2
timestamp 1734044400
transform 1 0 6984 0 1 1056
box -184 -128 1336 928
use JNWTR_CAPX1  xf ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1723932000
transform 1 0 0 0 1 4840
box 0 0 1080 1080
use JNWTR_CAPX1  xg1
timestamp 1723932000
transform 1 0 1760 0 1 4840
box 0 0 1080 1080
use JNWATR_NCH_4C5F0  xg2
timestamp 1734044400
transform 1 0 1760 0 1 5920
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xg3
timestamp 1734044400
transform 1 0 1760 0 1 6976
box -184 -128 1336 928
<< labels >>
flabel metal1 3700 7044 3878 7264 0 FreeSans 160 0 0 0 VDD
flabel metal1 7466 -328 7568 -214 0 FreeSans 160 0 0 0 V_pluss
flabel metal1 4712 1018 4852 1156 0 FreeSans 160 0 0 0 V_minus
flabel metal1 756 6752 904 6868 0 FreeSans 160 0 0 0 Diff_Out
flabel metal1 1696 -424 1734 -364 0 FreeSans 160 0 0 0 VSS
<< properties >>
string FIXED_BBOX 0 0 8136 7520
<< end >>
